// Code your design here

// for test
module adder;
  
  
endmodule: adder
//
