// Code your testbench here
// or browse Examples

// just test

class tb.c extends uvm_test_top
  
endclass: tb.c

//
